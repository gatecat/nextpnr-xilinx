`timescale 1 ps / 1 ps

(* blackbox *)
module zynq_ultra_ps_e_0 (
	output pl_clk0,
	input maxihpm0_fpd_aclk,
	input maxihpm1_fpd_aclk,
	input maxigp0_arready,
	input maxigp0_awready,
	input maxigp0_bid,
	input maxigp0_bresp,
	input maxigp0_bvalid,
	input maxigp0_rdata,
	input maxigp0_rid,
	input maxigp0_rlast,
	input maxigp0_rresp,
	input maxigp0_rvalid,
	input maxigp0_wready,
	input maxigp1_arready,
	input maxigp1_awready,
	input maxigp1_bid,
	input maxigp1_bresp,
	input maxigp1_bvalid,
	input maxigp1_rdata,
	input maxigp1_rid,
	input maxigp1_rlast,
	input maxigp1_rresp,
	input maxigp1_rvalid,
	input maxigp1_wready,
	input pl_ps_irq0
);
endmodule
